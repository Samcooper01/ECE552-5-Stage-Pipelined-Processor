/*
   CS/ECE 552 Spring '22
  
   Filename        : execute.v
   Description     : This is the overall module for the execute stage of the processor.
*/
module execute (clk, rst,
                BSrc, BSel, Cin, InvA, InvB, ALUOp, // control signal inputs
                opcode, read_data_1, read_data_2, instruction_lower_5_ext, instruction_lower_8_ext, instruction_lower_8, // data inputs
                ImmJmp, ALU_output, ALU_input_2, SLBI_concat); // data outputs

   // Inputs:
   input wire clk;
   input wire rst;
   input wire [1:0] BSrc;     // control signal 
   input wire BSel;     // control signal
   input wire Cin;      // control signal
   input wire InvA;     // control signal
   input wire InvB;     // control signal
   input wire [3:0] ALUOp;    // control signal for the ALU itself generated by ALU operation block
   input wire [4:0] opcode;                     // the opcode from the instruction
   input wire [15:0] read_data_1;               // read data 1 from reg file to ALU input 1
   input wire [15:0] read_data_2;               // read data 2 from reg file to mux ALU input 2
   input wire [15:0] instruction_lower_5_ext;   // lower 5 bits for mux ALU input 2
   input wire [15:0] instruction_lower_8_ext;   // lower 8 bits for mux ALU input 2
   input wire [7:0] instruction_lower_8;        // lower 8 bits of instruction for SLBI concat block
   
   // Outputs:
   output wire ImmJmp;               // control signal from branch conditional block from ALU flags
   output wire [15:0] ALU_output;    // output of the ALU
   output wire [15:0] ALU_input_2;   // input 2 of the ALU for write data in data memory
   output wire [15:0] SLBI_concat;   // result of SLBI instruction for ConstSel mux

   // Internal wires:
   wire [15:0] BSel_const_mux;       // output of the BSel mux
   wire SF;                          // sign flag
   wire ZF;                          // zero flag
   wire OF;                          // overflow flag
   wire CF;                          // carry flag

   // localparams
   localparam [15:0] zero = 16'b0;    // 0 value for BSel mux
   localparam [15:0] eight = 4'h8; // 8 value for BSel mux
   
   // instantiate ALU
   ALU iALU(.A(read_data_1), .B(ALU_input_2), .invA(InvA), .invB(InvB), .c_in(Cin), .SF(SF), .ZF(ZF), .OF(OF), .CF(CF), .ALU_mode(ALUOp), .out(ALU_output));

   // BSel mux to produce the fourth choice input for ALU input B
   assign BSel_const_mux = (BSel) ? eight : zero;

   // BSrc mux to select the input for ALU input B
   assign ALU_input_2 = (BSrc == 2'b00) ? read_data_2 :
                        (BSrc == 2'b01) ? instruction_lower_5_ext :
                        (BSrc == 2'b10) ? instruction_lower_8_ext :
                        (BSel_const_mux); // we default to the BSel mux for BSrc == 2'b11

   // TODO: create the BrchCnd block
   branchCnd ibranchCnd(.opcode(opcode), .SF(SF), .ZF(ZF), .OF(OF), .CF(CF), .immJump(ImmJmp));

   // custom hardware for SLBI instruction to produce SLBI_concat signal
   assign SLBI_concat = {ALU_output[15:8], instruction_lower_8};

endmodule
